-- In this VHDL file, AND, OR, NAND, NOR, XOR, XNOR and NOT gates 
--are implemented with the required delay. 

--AND GATE WITH 2 INPUTS
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY and2 IS
	PORT ( a, b: IN STD_LOGIC;
			  c: OUT STD_LOGIC);
END ENTITY and2;

ARCHITECTURE delayed OF and2 IS
BEGIN
	c <= a AND b AFTER 6 NS;
END ARCHITECTURE delayed;	

--AND GATE WITH 3 INPUTS 

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY and3 IS
	PORT ( a, b, c: IN STD_LOGIC;
			     d: OUT STD_LOGIC);
END ENTITY and3;

ARCHITECTURE delayed OF and3 IS
BEGIN
	d <= a AND b AND c AFTER 6 NS;
END ARCHITECTURE delayed;	  

--OR GATE WITH 2 INPUTS

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY or2 IS
	PORT ( a, b: IN STD_LOGIC;
			  c: OUT STD_LOGIC);
END ENTITY or2;

ARCHITECTURE delayed OF or2 IS
BEGIN
	c <= a OR b AFTER 6 NS;
END ARCHITECTURE delayed;	

--OR GATE WITH 3 INPUTS	 

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY or3 IS
	PORT ( a, b, c: IN STD_LOGIC;
			     d: OUT STD_LOGIC);
END ENTITY or3;

ARCHITECTURE delayed OF or3 IS
BEGIN
	d <= a OR b OR c AFTER 6 NS;
END ARCHITECTURE delayed;	

--OR GATE WITH 4 INPUTS	 

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY or4 IS
	PORT ( a, b, c, d: IN STD_LOGIC;
			        e: OUT STD_LOGIC);
END ENTITY or4;

ARCHITECTURE delayed OF or4 IS
BEGIN
	e <= a OR b OR c OR d AFTER 6 NS;
END ARCHITECTURE delayed;  

--OR GATE WITH 5 INPUTS	 

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY or5 IS
	PORT ( a, b, c, d, e: IN STD_LOGIC;
			        f: OUT STD_LOGIC);
END ENTITY or5;

ARCHITECTURE delayed OF or5 IS
BEGIN
	f <= a OR b OR c OR d OR e AFTER 6 NS;
END ARCHITECTURE delayed;  

--NAND GATE WITH 2 INPUTS

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY nand2 IS
	PORT ( a, b: IN STD_LOGIC;
			  c: OUT STD_LOGIC);
END ENTITY nand2;

ARCHITECTURE delayed OF nand2 IS
BEGIN
	c <= a NAND b AFTER 4 NS;
END ARCHITECTURE delayed; 

--NAND GATE WITH 3 INPUTS

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY nand3 IS
	PORT ( a, b, c: IN STD_LOGIC;
			  d: OUT STD_LOGIC);
END ENTITY nand3;

ARCHITECTURE delayed OF nand3 IS
BEGIN
	d <= (a NAND b) NAND c AFTER 4 NS;
END ARCHITECTURE delayed;  

--NAND GATE WITH 4 INPUTS

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY nand4 IS
	PORT ( a, b, c, d: IN STD_LOGIC;
			  y: OUT STD_LOGIC);
END ENTITY nand4;
--ASK THE DOCTOR
ARCHITECTURE delayed OF nand4 IS
BEGIN
	y <= (a NAND b) NAND (c NAND d) AFTER 4 NS;
END ARCHITECTURE delayed;  

--NOR GATE WITH 2 INPUTS

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY nor2 IS
	PORT ( a, b: IN STD_LOGIC;
			  c: OUT STD_LOGIC);
END ENTITY nor2;

ARCHITECTURE delayed OF nor2 IS
BEGIN
	c <= a NOR b AFTER 4 NS;
END ARCHITECTURE delayed; 

--XOR GATE WITH 2 INPUTS

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY xor2 IS
	PORT ( a, b: IN STD_LOGIC;
			  c: OUT STD_LOGIC);
END ENTITY xor2;

ARCHITECTURE delayed OF xor2 IS
BEGIN
	c <= a XOR b AFTER 8 NS;
END ARCHITECTURE delayed;  

--XOR GATE WITH 3 INPUTS	 

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY xor3 IS
	PORT ( a, b, c: IN STD_LOGIC;
			     d: OUT STD_LOGIC);
END ENTITY xor3;

ARCHITECTURE delayed OF xor3 IS
BEGIN
	d <= a XOR b XOR c AFTER 6 NS;
END ARCHITECTURE delayed;

--XNOR GATE WITH 2 INPUTS

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY xnor2 IS
	PORT ( a, b: IN STD_LOGIC;
			  c: OUT STD_LOGIC);
END ENTITY xnor2;

ARCHITECTURE delayed OF xnor2 IS
BEGIN
	c <= a XNOR b AFTER 7 NS;
END ARCHITECTURE delayed;  

--NOT GATE 

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY not1 IS
	PORT ( a: IN STD_LOGIC;
		   b: OUT STD_LOGIC);
END ENTITY not1;

ARCHITECTURE delayed OF not1 IS
BEGIN
	b <= NOT a AFTER 3 NS;
END ARCHITECTURE delayed;


